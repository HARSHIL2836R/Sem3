module karatsuba_16 (X, Y, Z);
input [15:0] X,Y;
output [31:0] Z;


endmodule
